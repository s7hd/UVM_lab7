package yapp_pkg;
  import uvm_pkg::*;
  //declaration 
  typedef uvm_config_db#(virtual yapp_if) yapp_vif_config;

  `include "uvm_macros.svh"
  
  `include "../task1_integ/yapp_packet.sv"
  `include "../task1_integ/yapp_tx_monitor.sv"
  `include "../task1_integ/yapp_tx_sequencer.sv"
  `include "../task1_integ/yapp_tx_seqs.sv"
  `include "../task1_integ/yapp_tx_driver.sv"
  `include "../task1_integ/yapp_tx_agent.sv"
  `include "../task1_integ/yapp_tx_env.sv"
  
endpackage